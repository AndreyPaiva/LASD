module DecodificadorHexa7Seg(
input [3:0] in,
output[6:0] out
);
reg [6:0] hexa7seg;

always @(*)
	begin
		case(in[3:0])
			4'b0000	:	hexa7seg[6:0] = 7'b0000001;
			4'b0001	:	hexa7seg[6:0] = 7'b1001111;
			4'b0010	:	hexa7seg[6:0] = 7'b0010010;
			4'b0011	:	hexa7seg[6:0] = 7'b0000110;
			4'b0100	:	hexa7seg[6:0] = 7'b1001100;
			4'b0101	:	hexa7seg[6:0] = 7'b0100100;
			4'b0110	:	hexa7seg[6:0] = 7'b0100000;
			4'b0111	:	hexa7seg[6:0] = 7'b0001111;
			4'b1000	:	hexa7seg[6:0] = 7'b0000000;
			4'b1001	:	hexa7seg[6:0] = 7'b0000100;
			4'b1010	:	hexa7seg[6:0] = 7'b0001000;
			4'b1011	:	hexa7seg[6:0] = 7'b1100000;
			4'b1100	:	hexa7seg[6:0] = 7'b0110001;
			4'b1101	:	hexa7seg[6:0] = 7'b1000010;
			4'b1110	:	hexa7seg[6:0] = 7'b0110000;
			4'b1111	:	hexa7seg[6:0] = 7'b0111000;
			default	:  hexa7seg[6:0] = 7'b0000000;
		endcase
	end
	
	assign out[6:0] = hexa7seg[6:0];
	
endmodule